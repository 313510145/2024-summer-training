module top_809960632_810038711_1598227639_893650103 (n51, n12, n67, n78, n22, n80, n72, n75, n2, n18, n57, n34, n4, n35, n56);
input n51, n12, n67, n78, n22, n80, n72, n75, n2, n18, n57, n34, n4, n35;
output n56;
wire n8, n60, n37, n5, n45, n54, n88, n43, n20, n53, n58, n41, n83, n29, n40, n27, n16, n10, n15, n69, n0, n66, n85, n24, n87, n26, n50, n28, n17, n36, n23, n89, n61, n7, n84, n76, n62, n30, n11, n46, n71, n31, n44, n55, n52, n64, n13, n19, n79, n39, n81, n1, n70, n47, n82, n90, n14, n21, n59, n25, n49, n3, n38, n74, n42, n6, n65, n9;
and_6 g54 (n8, n89, n56);
and_6 g73 (n6, n42, n8);
xnor_4 g28 (n60, n5, n6);
or_6 g22 (n37, n12, n60);
not_8 g40 (n51, n37);
xnor_4 g1 (n45, n53, n5);
and_6 g31 (n54, n43, n45);
or_6 g57 (n88, n78, n54);
not_8 g24 (n67, n88);
and_6 g19 (n22, n20, n43);
or_6 g12 (n80, n67, n20);
or_6 g66 (n58, n41, n53);
and_6 g8 (n72, n67, n58);
or_6 g56 (n22, n83, n41);
nor_5 g68 (n29, n67, n83);
not_8 g33 (n75, n29);
xor_4 g37 (n40, n69, n42);
nor_5 g3 (n12, n27, n40);
and_6 g20 (n53, n16, n27);
not_8 g4 (n10, n16);
and_6 g44 (n51, n15, n10);
not_8 g16 (n45, n15);
xnor_4 g17 (n0, n50, n69);
not_8 g69 (n66, n0);
and_6 g65 (n85, n87, n66);
or_6 g67 (n24, n78, n85);
not_8 g9 (n2, n24);
and_6 g25 (n18, n26, n87);
or_6 g7 (n80, n2, n26);
and_6 g15 (n28, n36, n50);
or_6 g76 (n17, n24, n28);
not_8 g58 (n72, n17);
nor_5 g48 (n18, n23, n36);
nor_5 g62 (n29, n2, n23);
and_6 g39 (n9, n65, n89);
xor_4 g2 (n61, n30, n9);
nor_5 g45 (n12, n7, n61);
nor_5 g13 (n84, n76, n7);
and_6 g74 (n0, n10, n84);
or_6 g64 (n50, n62, n76);
nor_5 g72 (n53, n66, n62);
xnor_4 g55 (n11, n55, n30);
and_6 g61 (n46, n31, n11);
or_6 g49 (n71, n78, n46);
not_8 g27 (n57, n71);
and_6 g6 (n34, n44, n31);
or_6 g63 (n80, n57, n44);
or_6 g32 (n52, n64, n55);
and_6 g14 (n72, n57, n52);
or_6 g75 (n34, n13, n64);
nor_5 g52 (n29, n57, n13);
xor_4 g38 (n19, n82, n65);
nor_5 g59 (n12, n79, n19);
and_6 g11 (n39, n1, n79);
or_6 g51 (n11, n81, n39);
not_8 g5 (n84, n81);
and_6 g23 (n55, n70, n1);
or_6 g47 (n11, n47, n70);
not_8 g70 (n76, n47);
xor_4 g53 (n90, n49, n82);
and_6 g41 (n14, n59, n90);
or_6 g10 (n21, n78, n14);
not_8 g21 (n4, n21);
and_6 g30 (n35, n25, n59);
or_6 g42 (n80, n4, n25);
and_6 g43 (n3, n38, n49);
nand_5 g18 (n72, n4, n3);
nor_5 g60 (n35, n74, n38);
nor_5 g34 (n29, n4, n74);
endmodule
