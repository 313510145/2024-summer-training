module top_809960632_810038711_1598227639_893650103 (n4, n78, n35, n80, n57, n34, n2, n18, n67, n22, n77);
input n4, n78, n35, n80, n57, n34, n2, n18, n67, n22;
output n77;
wire n86, n90, n14, n21, n59, n25, n11, n46, n71, n31, n44, n73, n66, n85, n24, n87, n26, n45, n54, n88, n43, n20;
or_6 g0 (n86, n73, n77);
or_6 g35 (n90, n11, n86);
and_6 g41 (n14, n59, n90);
or_6 g10 (n21, n78, n14);
not_8 g21 (n4, n21);
and_6 g30 (n35, n25, n59);
or_6 g42 (n80, n4, n25);
and_6 g61 (n46, n31, n11);
or_6 g49 (n71, n78, n46);
not_8 g27 (n57, n71);
and_6 g6 (n34, n44, n31);
or_6 g63 (n80, n57, n44);
or_6 g36 (n66, n45, n73);
and_6 g65 (n85, n87, n66);
or_6 g67 (n24, n78, n85);
not_8 g9 (n2, n24);
and_6 g25 (n18, n26, n87);
or_6 g7 (n80, n2, n26);
and_6 g31 (n54, n43, n45);
or_6 g57 (n88, n78, n54);
not_8 g24 (n67, n88);
and_6 g19 (n22, n20, n43);
or_6 g12 (n80, n67, n20);
endmodule
